$date
	Mon Nov 17 16:12:27 2025
$end
$version
	Icarus Verilog
$end
$timescale
	1ps
$end
$scope module dmem_tb $end
$var wire 32 ! rdata [31:0] $end
$var reg 1 " MemRead $end
$var reg 1 # MemWrite $end
$var reg 32 $ addr [31:0] $end
$var reg 1 % clk $end
$var reg 32 & wdata [31:0] $end
$scope module UUT $end
$var wire 1 " MemRead $end
$var wire 1 # MemWrite $end
$var wire 32 ' addr [31:0] $end
$var wire 1 % clk $end
$var wire 32 ( wdata [31:0] $end
$var wire 32 ) rdata [31:0] $end
$upscope $end
$upscope $end
$enddefinitions $end
$comment Show the parameter values. $end
$dumpall
$end
#0
$dumpvars
b0 )
b0 (
b0 '
b0 &
0%
b0 $
0#
0"
b0 !
$end
#5000
1%
#10000
b11011110101011011011111011101111 !
b11011110101011011011111011101111 )
0%
1"
#15000
1%
#20000
b0 !
b0 )
0%
b10010001101000101011001111000 &
b10010001101000101011001111000 (
b1000 $
b1000 '
1#
0"
#25000
1%
#30000
b10010001101000101011001111000 !
b10010001101000101011001111000 )
0%
1"
0#
#35000
1%
#40000
0%
